// ----  Probes  ----
`define PROBE_F_PC if_pc
`define PROBE_F_INSN if_insn

`define PROBE_D_PC id_pc
`define PROBE_D_OPCODE id_opcode
`define PROBE_D_RD id_rd
`define PROBE_D_FUNCT3 id_funct3
`define PROBE_D_RS1 id_rs1
`define PROBE_D_RS2 id_rs2
`define PROBE_D_FUNCT7 id_funct7
`define PROBE_D_IMM id_imm
`define PROBE_D_SHAMT id_shamt
// ----  Probes  ----

// ----  Top module  ----
`define TOP_MODULE  pd2
// ----  Top module  ----
